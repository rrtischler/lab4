module InstFetch(NPC, IR, MEM_ADDR, MEM_CLK, RST, CLK, ULA, COND, MEM_OUT);

	output reg [15:0] NPC;
	output reg [31:0] IR;
	output [15:0] MEM_ADDR;
	output MEM_CLK;
	
	input RST;
	input CLK;
	input [15:0] ULA;
	input COND;
	input [31:0] MEM_OUT;
	
	
	
	
	
	
endmodule
