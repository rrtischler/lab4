module WriteBack()



endmodule
