module MemAcc();


endmodule
