module Exec( );



endmodule
